-- cell_ctrl.vhd
-- Autori: Jakub Cabal
-- Posledni zmena: 12.12.2014
-- Popis: Obvod pro rizeni zobrazovani pole
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity CELL_CTRL is
   Port (
      CLK         : in  STD_LOGIC;
      PIXEL_X     : in  STD_LOGIC_VECTOR (9 downto 0);
      PIXEL_Y     : in  STD_LOGIC_VECTOR (9 downto 0);
      KURZOR_ADDR : in  STD_LOGIC_VECTOR (7 downto 0);
      KURZOR      : out STD_LOGIC;
      PIXEL_SET_X : out STD_LOGIC;
      PIXEL_SET_Y : out STD_LOGIC;
      KOMP_SET_X  : out STD_LOGIC;
      KOMP_SET_Y  : out STD_LOGIC;
      KOMP_ON     : out STD_LOGIC;
      ADDR        : out STD_LOGIC_VECTOR (7 downto 0);
      KOMP0       : in  STD_LOGIC_VECTOR (5 downto 0);
      KOMP1       : in  STD_LOGIC_VECTOR (5 downto 0);
      KOMP2       : in  STD_LOGIC_VECTOR (5 downto 0);
      KOMP3       : in  STD_LOGIC_VECTOR (5 downto 0);
      KOMP4       : in  STD_LOGIC_VECTOR (5 downto 0);
      KOMP_OUT    : out STD_LOGIC_VECTOR (5 downto 0);
      MAIN_SC     : in  STD_LOGIC;
      GAME_SC     : in  STD_LOGIC;
      LVL2_SC     : in  STD_LOGIC;
      LVL3_SC     : in  STD_LOGIC;
      LVL4_SC     : in  STD_LOGIC;
      WIN_SC      : in  STD_LOGIC;
      LOSE_SC     : in  STD_LOGIC
   );                    
end CELL_CTRL;

architecture FULL of CELL_CTRL is

   signal pix_x           : STD_LOGIC_VECTOR(9 downto 0);
   signal pix_y           : STD_LOGIC_VECTOR(9 downto 0);
   
   signal addr_x          : STD_LOGIC_VECTOR(3 downto 0);
   signal addr_y          : STD_LOGIC_VECTOR(3 downto 0);
   signal addr_x2         : STD_LOGIC_VECTOR(3 downto 0) := (others => '0');
   signal addr_y2         : STD_LOGIC_VECTOR(3 downto 0) := (others => '0');

   signal obj_addr_x      : STD_LOGIC_VECTOR(4 downto 0);
   signal obj_addr_x2     : STD_LOGIC_VECTOR(4 downto 0) := (others => '0');

   signal obj_addr_y      : STD_LOGIC_VECTOR(3 downto 0);
   signal obj_addr_y2     : STD_LOGIC_VECTOR(3 downto 0) := (others => '0');
   
   signal pix_set_x       : STD_LOGIC;
   signal pix_set_y       : STD_LOGIC;

   signal sig_kurzor_x    : STD_LOGIC_VECTOR(3 downto 0);
   signal sig_kurzor_y    : STD_LOGIC_VECTOR(3 downto 0);
   signal kurzor_set_x    : STD_LOGIC;
   signal kurzor_set_y    : STD_LOGIC;

   signal k_set_x         : STD_LOGIC;
   signal k_set_y         : STD_LOGIC;

   signal sig_kset_x      : STD_LOGIC;
   signal sig_kset_y      : STD_LOGIC;

   signal sig_komp_on     : STD_LOGIC;
   signal pre_komp_out    : STD_LOGIC_VECTOR(5 downto 0);
   signal rom_addr        : STD_LOGIC_VECTOR(11 downto 0);
   signal rom_data        : STD_LOGIC_VECTOR(8 downto 0);
   signal game_screens    : STD_LOGIC_VECTOR(2 downto 0);

   -- Blokova pamet -- konfigurace obrazovek
   type rom_type is array (0 to 4095) of STD_LOGIC_VECTOR(0 to 8);
   constant ROM : rom_type :=
   (
      -- main screen
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --1.r

      "000000000",
      "000000000",
      "000000000",
      "110010100",
      "000001100",
      "000010100",
      "000000000",
      "000011100", 
      "000000000",
      "110010100", 
      "000001100", 
      "000010100",
      "000000000",
      "000011100", 
      "000001100", 
      "000010100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --2.r

      "000000000",
      "000000000",
      "000000000",
      "010001100", 
      "000000000",
      "010001100", 
      "000000000",
      "010001100", 
      "000000000",
      "010001100", 
      "000000000",
      "010001100", 
      "000000000",
      "010001100", 
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --3.r

      "000000000",
      "000000000",
      "000000000",
      "000011100", 
      "000001100", 
      "010010100", 
      "000000000",
      "010001100", 
      "000000000",
      "000011100", 
      "000001100", 
      "010010100", 
      "000000000",
      "000011100", 
      "000001100", 
      "000000000",
      "000000000", 
      "000000000", 
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --4.r

      "000000000",
      "000000000",
      "000000000",
      "010001100", 
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --5.r

      "000000000",
      "000000000",
      "000000000",
      "010001100", 
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000011100",
      "000001100",
      "010010100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --6.r

      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --7.r

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --8.r

      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000011100",
      "000000000",
      "000000000",
      "000001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --9.r

      "000011100",
      "000010100",
      "000000000",
      "110010100", 
      "000011100",
      "000000000",
      "110010100",
      "000000000",
      "000010100", 
      "000000000",
      "000011100",
      "000010100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "110010100",
      "000000000",
      "000010100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --10.r

      "010001100",
      "000000000",
      "000001100", 
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "100010100", 
      "000011100", 
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --11.r

      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000011100",
      "000001100",
      "000011100",
      "000000000", 
      "010001100",
      "000000000",
      "000000000", 
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000011100",
      "000001100",
      "000011100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --12.r

      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --13.r

      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --14.r

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001001100",
      "001101100",
      "001110100",
      "001111100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --15.r

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --16.r

      --game screen

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --1.r

      "000000000",
      "000110100",
      "000111100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --2.r

      "000000000",
      "000101100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000101", -- KOMP0
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --3.r

      "000000000",
      "000101100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --4.r

      "000000000",
      "000101100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000110", -- KOMP1
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --5.r

      "000000000",
      "000101100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --6.r

      "000000000",
      "000101100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000111", -- KOMP2
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --7.r

      "000000000",
      "000101100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --8.r

      "000000000",
      "000101100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000001", -- KOMP3
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --9.r

      "000000000",
      "000101100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --10.r

      "000000000",
      "000100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000010", -- KOMP4
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --11.r

      "001011100",
      "001010100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --12.r

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --13.r

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001000100",
      "000111100",
      "000111100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --14.r

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --15.r

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --16.r
      -- win screen
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --1.ř.

      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --2.ř.

      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "110010100",
      "000001100",
      "000010100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --3.ř.

      "000000000",
      "000000000",
      "100010100",
      "000011100",
      "010010100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --4.ř.

      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "100010100",
      "000001100",
      "000011100",
      "000001100",
      "010010100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --5.ř.

      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000001100",
      "000000000",
      "000000000",
      "000000000",
      "000001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --6.ř.

      "000000000",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --7.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --8.ř.

      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000011100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "110010100",
      "000001100",
      "000011100",
      "000001100",
      "000010100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --9.ř.

      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000011100",
      "000010100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --10.ř.

      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "100010100",
      "000011100",
      "000000000",
      "100010100",
      "000001100",
      "010010100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --11.ř.

      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --12.ř.

      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "110010100",
      "000010100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --13.ř.

      "000000000",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "000000000",
      "100010100",
      "000011100",
      "000001100",
      "010010100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --14.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --15.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000", --16.r
      -- lose screen
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000011100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --1.ř.

      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --2.ř.

      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "100010100",
      "010001100",
      "000010100",
      "110010100",
      "000001100",
      "000010100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --3.ř.

      "000000000",
      "000000000",
      "100010100",
      "000011100",
      "010010100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "100010100",
      "000001100",
      "010010100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --4.ř.

      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000001100",
      "000000000",
      "000000000",
      "110010100",
      "010010100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --5.ř.

      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000001100",
      "000000000",
      "000000000",
      "000000000",
      "000001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "110010100",
      "000001100",
      "010010100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --6.ř.

      "000000000",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "000000000",
      "000000000",
      "100010100",
      "000001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --7.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --8.ř.

      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000001100",
      "000000000",
      "000000000",
      "000000000",
      "000001100",
      "000001100",
      "000000000",
      "000011100",
      "000001100",
      "000010100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --9.ř.

      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --10.ř.

      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000001100",
      "000000000",
      "000000000",
      "000011100",
      "000001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --11.ř.

      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --12.ř.

      "000000000",
      "000000000",
      "000011100",
      "000001100",
      "010010100",
      "000000000",
      "000000000",
      "000001100",
      "000000000",
      "000000000",
      "000001100",
      "000001100",
      "000000000",
      "000000000",
      "000011100",
      "000001100",
      "010010100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --13.ř.

      "000000000",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --14.r.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --15.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --16.ř.
      -- lvl2
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --1.ř.

      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000011100",
      "000001100",
      "000010100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000011100",
      "000001100",
      "000010100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --2.ř.

      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --3.ř.

      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000011100",
      "000001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000011100",
      "000001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --4.ř.

      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --5.ř.

      "000011100",
      "000001100",
      "010010100",
      "000000000",
      "000011100",
      "000001100",
      "010010100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000011100",
      "000001100",
      "010010100",
      "000000000",
      "000011100",
      "000001100",
      "010010100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --6.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --7.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --8.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --9.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --10.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --11.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --12.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --13.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --14.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001001100",
      "001101100",
      "001110100",
      "001111100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --15.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --16.ř.
      -- lvl3
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --1.ř.

      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000011100",
      "000001100",
      "000010100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000011100",
      "000001100",
      "000010100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --2.ř.

      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --3.ř.

      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000011100",
      "000001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000011100",
      "000001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --4.ř.

      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --5.ř.

      "000011100",
      "000001100",
      "010010100",
      "000000000",
      "000011100",
      "000001100",
      "010010100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000011100",
      "000001100",
      "010010100",
      "000000000",
      "000011100",
      "000001100",
      "010010100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --6.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --7.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --8.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --9.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --10.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --11.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --12.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --13.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --14.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001001100",
      "001101100",
      "001110100",
      "001111100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --15.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --16.ř.
      -- lvl4
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --1.ř.

      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000011100",
      "000001100",
      "000010100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000011100",
      "000001100",
      "000010100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --2.ř.

      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --3.ř.

      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000011100",
      "000001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "010001100",
      "000000000",
      "000011100",
      "000001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --4.ř.

      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --5.ř.

      "000011100",
      "000001100",
      "010010100",
      "000000000",
      "000011100",
      "000001100",
      "010010100",
      "000000000",
      "000000000",
      "010001100",
      "000000000",
      "000000000",
      "000011100",
      "000001100",
      "010010100",
      "000000000",
      "000011100",
      "000001100",
      "010010100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --6.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --7.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --8.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --9.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --10.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "000000000",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --11.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "000000000",
      "000000000",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --12.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --13.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001100100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --14.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "001001100",
      "001101100",
      "001110100",
      "001111100",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --15.ř.

      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",
      "000000000",   --16.ř.
      others => (others => '0')
   );

begin

   pix_x <= PIXEL_X;
   pix_y <= PIXEL_Y;

   ------------------------------------------------------------------
   -- ZOBRAZOVANI HERNIHO POLE
   ------------------------------------------------------------------
   
   process (CLK)
   begin
      if rising_edge(CLK) then
         if (pix_x = 0) then
            pix_set_x <= '0';
            k_set_x   <= '1';
            addr_x <= (others => '0');
            obj_addr_x <= std_logic_vector(to_unsigned(0, 5));
         elsif (pix_x = 32) then
            pix_set_x <= '0';
            k_set_x   <= '1';
            addr_x <= (others => '0');
            obj_addr_x <= std_logic_vector(to_unsigned(1, 5));
         elsif (pix_x = 64) then
            pix_set_x <= '0';
            k_set_x   <= '1';
            addr_x <= (others => '0');
            obj_addr_x <= std_logic_vector(to_unsigned(2, 5));
         elsif (pix_x = 96) then
            pix_set_x <= '1';
            k_set_x   <= '1';
            addr_x <= std_logic_vector(to_unsigned(0, 4));
            obj_addr_x <= std_logic_vector(to_unsigned(3, 5));
         elsif (pix_x = 128) then
            pix_set_x <= '1';
            k_set_x   <= '1';
            addr_x <= std_logic_vector(to_unsigned(1, 4));
            obj_addr_x <= std_logic_vector(to_unsigned(4, 5));
         elsif (pix_x = 160) then
            pix_set_x <= '1';
            k_set_x   <= '1';
            addr_x <= std_logic_vector(to_unsigned(2, 4));
            obj_addr_x <= std_logic_vector(to_unsigned(5, 5));
         elsif (pix_x = 192) then
            pix_set_x <= '1';
            k_set_x   <= '1';
            addr_x <= std_logic_vector(to_unsigned(3, 4));
            obj_addr_x <= std_logic_vector(to_unsigned(6, 5));
         elsif (pix_x = 224) then
            pix_set_x <= '1';
            k_set_x   <= '1';
            addr_x <= std_logic_vector(to_unsigned(4, 4));
            obj_addr_x <= std_logic_vector(to_unsigned(7, 5));
         elsif (pix_x = 256) then
            pix_set_x <= '1';
            k_set_x   <= '1';
            addr_x <= std_logic_vector(to_unsigned(5, 4));
            obj_addr_x <= std_logic_vector(to_unsigned(8, 5));
         elsif (pix_x = 288) then
            pix_set_x <= '1';
            k_set_x   <= '1';
            addr_x <= std_logic_vector(to_unsigned(6, 4));
            obj_addr_x <= std_logic_vector(to_unsigned(9, 5));
         elsif (pix_x = 320) then
            pix_set_x <= '1';
            k_set_x   <= '1';
            addr_x <= std_logic_vector(to_unsigned(7, 4));
            obj_addr_x <= std_logic_vector(to_unsigned(10, 5));
         elsif (pix_x = 352) then
            pix_set_x <= '1';
            k_set_x   <= '1';
            addr_x <= std_logic_vector(to_unsigned(8, 4));
            obj_addr_x <= std_logic_vector(to_unsigned(11, 5));
         elsif (pix_x = 384) then
            pix_set_x <= '1';
            k_set_x   <= '1';
            addr_x <= std_logic_vector(to_unsigned(9, 4));
            obj_addr_x <= std_logic_vector(to_unsigned(12, 5));
         elsif (pix_x = 416) then
            pix_set_x <= '1';
            k_set_x   <= '1';
            addr_x <= std_logic_vector(to_unsigned(10, 4));
            obj_addr_x <= std_logic_vector(to_unsigned(13, 5));
         elsif (pix_x = 448) then
            pix_set_x <= '1';
            k_set_x   <= '1';
            addr_x <= std_logic_vector(to_unsigned(11, 4));
            obj_addr_x <= std_logic_vector(to_unsigned(14, 5));
         elsif (pix_x = 480) then
            pix_set_x <= '1';
            k_set_x   <= '1';
            addr_x <= std_logic_vector(to_unsigned(12, 4));
            obj_addr_x <= std_logic_vector(to_unsigned(15, 5));
         elsif (pix_x = 512) then
            pix_set_x <= '1';
            k_set_x   <= '1';
            addr_x <= std_logic_vector(to_unsigned(13, 4));
            obj_addr_x <= std_logic_vector(to_unsigned(16, 5));
         elsif (pix_x = 544) then
            pix_set_x <= '0';
            k_set_x   <= '1';
            addr_x <= (others => '0');
            obj_addr_x <= std_logic_vector(to_unsigned(17, 5));
         elsif (pix_x = 576) then
            pix_set_x <= '0';
            k_set_x   <= '1';
            addr_x <= (others => '0');
            obj_addr_x <= std_logic_vector(to_unsigned(18, 5));
         elsif (pix_x = 608) then
            pix_set_x <= '0';
            k_set_x   <= '1';
            addr_x <= (others => '0');
            obj_addr_x <= std_logic_vector(to_unsigned(19, 5));
         else
            pix_set_x <= '0';
            k_set_x   <= '0';
            addr_x <= (others => '0');
            obj_addr_x <= (others => '0');
         end if;
      end if;
   end process;
   
   process (CLK)
   begin
      if rising_edge(CLK) then
         if (pix_y = 0) then
            pix_set_y <= '0';
            k_set_y <= '1';
            addr_y <= (others => '0');
            obj_addr_y <= std_logic_vector(to_unsigned(0, 4));
         elsif (pix_y = 32) then
            pix_set_y <= '1';
            k_set_y <= '1';
            addr_y <= std_logic_vector(to_unsigned(0, 4));
            obj_addr_y <= std_logic_vector(to_unsigned(1, 4));
         elsif (pix_y = 64) then
            pix_set_y <= '1';
            k_set_y <= '1';
            addr_y <= std_logic_vector(to_unsigned(1, 4));
            obj_addr_y <= std_logic_vector(to_unsigned(2, 4));
         elsif (pix_y = 96) then
            pix_set_y <= '1';
            k_set_y <= '1';
            addr_y <= std_logic_vector(to_unsigned(2, 4));
            obj_addr_y <= std_logic_vector(to_unsigned(3, 4));
         elsif (pix_y = 128) then
            pix_set_y <= '1';
            k_set_y <= '1';
            addr_y <= std_logic_vector(to_unsigned(3, 4));
            obj_addr_y <= std_logic_vector(to_unsigned(4, 4));
         elsif (pix_y = 160) then
            pix_set_y <= '1';
            k_set_y <= '1';
            addr_y <= std_logic_vector(to_unsigned(4, 4));
            obj_addr_y <= std_logic_vector(to_unsigned(5, 4));
         elsif (pix_y = 192) then
            pix_set_y <= '1';
            k_set_y <= '1';
            addr_y <= std_logic_vector(to_unsigned(5, 4));
            obj_addr_y <= std_logic_vector(to_unsigned(6, 4));
         elsif (pix_y = 224) then
            pix_set_y <= '1';
            k_set_y <= '1';
            addr_y <= std_logic_vector(to_unsigned(6, 4));
            obj_addr_y <= std_logic_vector(to_unsigned(7, 4));
         elsif (pix_y = 256) then
            pix_set_y <= '1';
            k_set_y <= '1';
            addr_y <= std_logic_vector(to_unsigned(7, 4));
            obj_addr_y <= std_logic_vector(to_unsigned(8, 4));
         elsif (pix_y = 288) then
            pix_set_y <= '1';
            k_set_y <= '1';
            addr_y <= std_logic_vector(to_unsigned(8, 4));
            obj_addr_y <= std_logic_vector(to_unsigned(9, 4));
         elsif (pix_y = 320) then
            pix_set_y <= '1';
            k_set_y <= '1';
            addr_y <= std_logic_vector(to_unsigned(9, 4));
            obj_addr_y <= std_logic_vector(to_unsigned(10, 4));
         elsif (pix_y = 352) then
            pix_set_y <= '1';
            k_set_y <= '1';
            addr_y <= std_logic_vector(to_unsigned(10, 4));
            obj_addr_y <= std_logic_vector(to_unsigned(11, 4));
         elsif (pix_y = 384) then
            pix_set_y <= '1';
            k_set_y <= '1';
            addr_y <= std_logic_vector(to_unsigned(11, 4));
            obj_addr_y <= std_logic_vector(to_unsigned(12, 4));
         elsif (pix_y = 416) then
            pix_set_y <= '1';
            k_set_y <= '1';
            addr_y <= std_logic_vector(to_unsigned(12, 4));
            obj_addr_y <= std_logic_vector(to_unsigned(13, 4));
         elsif (pix_y = 448) then
            pix_set_y <= '0';
            k_set_y <= '1';
            addr_y <= (others => '0');
            obj_addr_y <= std_logic_vector(to_unsigned(14, 4));
         else
            pix_set_y <= '0';
            k_set_y <= '0';
            addr_y <= (others => '0');
            obj_addr_y <= (others => '0');
         end if;
      end if;
   end process;
   
   ADDR         <= addr_y2 & addr_x2;
   sig_kurzor_x <= KURZOR_ADDR(3 downto 0);
   sig_kurzor_y <= KURZOR_ADDR(7 downto 4);

   process (CLK)
   begin
      if rising_edge(CLK) then
         if (pix_set_x = '1') then
            addr_x2 <= addr_x;
         end if;
      end if;
   end process;

   process (CLK)
   begin
      if rising_edge(CLK) then
         if (pix_set_x = '1' AND pix_set_y = '1') then
            addr_y2 <= addr_y;
         end if;
      end if;
   end process;

   process (CLK)
   begin
      if rising_edge(CLK) then
         if (k_set_x = '1') then
            obj_addr_x2 <= obj_addr_x;
         end if;
      end if;
   end process;

   process (CLK)
   begin
      if rising_edge(CLK) then
         if (k_set_x = '1' AND k_set_y = '1') then
            obj_addr_y2 <= obj_addr_y;
         end if;
      end if;
   end process;

   process (CLK)
   begin
      if rising_edge(CLK) then
         PIXEL_SET_X  <= pix_set_x;  
         PIXEL_SET_Y  <= pix_set_x AND pix_set_y;
         sig_kset_x   <= k_set_x;
         sig_kset_y   <= k_set_x AND k_set_y;
         KOMP_SET_X   <= sig_kset_x;
         KOMP_SET_Y   <= sig_kset_y;
      end if;
   end process;

   process (CLK)
   begin
      if rising_edge(CLK) then
         if (pix_set_x = '1') then
            if (sig_kurzor_x = addr_x) then
               kurzor_set_x <= '1';
            else
               kurzor_set_x <= '0';
            end if;
         end if;
      end if;
   end process;

   process (CLK)
   begin
      if rising_edge(CLK) then
         if (pix_set_x = '1' AND pix_set_y = '1') then
            if (sig_kurzor_y = addr_y) then
               kurzor_set_y <= '1';
            else
               kurzor_set_y <= '0';
            end if;
         end if;
      end if;
   end process;

   KURZOR <= kurzor_set_x AND kurzor_set_y;

   --------------------------------------------------------------------
   -- ZOBRAZOVANI OBJEKTU MIMO HERNI POLE VCETNE MEZI HERNICH OBRAZOVEK
   --------------------------------------------------------------------

   KOMP_ON  <= sig_komp_on;

   process (MAIN_SC, GAME_SC, WIN_SC, LOSE_SC, LVL2_SC, LVL3_SC, LVL4_SC)
   begin
      if (MAIN_SC = '1') then
         game_screens <= "000"; -- uvodni obrazovka
      elsif(GAME_SC = '1') then
         game_screens <= "001"; -- herni obrazovka
      elsif(WIN_SC = '1') then
         game_screens <= "010"; -- vyherni obrazovka
      elsif(LOSE_SC = '1') then
         game_screens <= "011"; -- game over obrazovka
      elsif(LVL2_SC = '1') then
         game_screens <= "100"; -- lvl2 obrazovka
      elsif(LVL3_SC = '1') then
         game_screens <= "101"; -- lvl3 obrazovka
      elsif(LVL4_SC = '1') then
         game_screens <= "110"; -- lvl4 obrazovka
      else
         game_screens <= "000"; -- jinak uvodni obrazovka
      end if;
   end process;

   -- Nastaveni cteci pameti
   rom_addr <= game_screens & obj_addr_y2 & obj_addr_x2;

   -- Vycteni dat z pameti ROM
   process (CLK)
   begin
      if rising_edge(CLK) then
         rom_data <= ROM(to_integer(unsigned(rom_addr)));  
      end if;
   end process;

   pre_komp_out <= rom_data(8 downto 3);

   with rom_data(2 downto 0) select
   KOMP_OUT <= pre_komp_out when "100",
               KOMP0 when "101",
               KOMP1 when "110",
               KOMP2 when "111",
               KOMP3 when "001",
               KOMP4 when "010",
               "000000" when others;

   with rom_data(2 downto 0) select
   sig_komp_on <= '1' when "100",
                  '1' when "101",
                  '1' when "110",
                  '1' when "111",
                  '1' when "001",
                  '1' when "010",
                  '0' when others;

end FULL;