-- cell_generator.vhd
-- Autori: Jakub Cabal, Tomas Bannert
-- Posledni zmena: 04.12.2014
-- Popis: Generator grafickych policek
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity CELL_GENERATOR is
   Port (
      CLK            : in  STD_LOGIC;
      RST            : in  STD_LOGIC; 
      TYP_ROURY      : in  STD_LOGIC_VECTOR (3 downto 0);
      NATOCENI_ROURY : in  STD_LOGIC_VECTOR (1 downto 0);
      ROURA_VODA1    : in  STD_LOGIC_VECTOR (5 downto 0);
      ROURA_VODA2    : in  STD_LOGIC_VECTOR (5 downto 0);
      ZDROJ_VODY1    : in  STD_LOGIC_VECTOR (3 downto 0);
      ZDROJ_VODY2    : in  STD_LOGIC_VECTOR (3 downto 0);
      KURZOR         : in  STD_LOGIC;
      PIXEL_X2       : in  STD_LOGIC_VECTOR (9 downto 0);
      PIXEL_Y2       : in  STD_LOGIC_VECTOR (9 downto 0);
      PIXEL_SET_X    : in  STD_LOGIC;
      PIXEL_SET_Y    : in  STD_LOGIC;
      KOMP_SET_X     : in  STD_LOGIC;
      KOMP_SET_Y     : in  STD_LOGIC;
      KOMP_ON        : in  STD_LOGIC;
      KOMP_IN        : in  STD_LOGIC_VECTOR (5 downto 0);
      GAME_ON        : in  STD_LOGIC;
      LOAD_WATER     : in  STD_LOGIC_VECTOR (7 downto 0);
      RGB            : out STD_LOGIC_VECTOR (2 downto 0)
   );                    
end CELL_GENERATOR;

architecture FULL of CELL_GENERATOR is

   signal cell_x_l   : unsigned(9 downto 0);
   signal cell_x_r   : unsigned(9 downto 0);
   signal cell_y_t   : unsigned(9 downto 0);
   signal cell_y_b   : unsigned(9 downto 0);
   signal rom_addr   : unsigned(8 downto 0);
   signal img_row    : unsigned(4 downto 0);
   signal img_col    : unsigned(4 downto 0);
   signal sig_komp_in        : STD_LOGIC_VECTOR(5 downto 0);
   signal rom_data           : STD_LOGIC_VECTOR(31 downto 0);
   signal rom_bit            : STD_LOGIC;
   signal sq_cell_on         : STD_LOGIC;
   signal sig_kurzor         : STD_LOGIC;
   signal sig_komp_on        : STD_LOGIC;
   signal pix_x              : unsigned(9 downto 0);
   signal pix_y              : unsigned(9 downto 0);
   signal pix_x2             : unsigned(9 downto 0);
   signal pix_y2             : unsigned(9 downto 0);
   signal sig_typ_roury      : STD_LOGIC_VECTOR(3 downto 0);
   signal sig_typ_roury2     : STD_LOGIC_VECTOR(3 downto 0);
   signal sig_natoceni_roury : STD_LOGIC_VECTOR(1 downto 0);
   signal load_water_lenght  : unsigned(9 downto 0);
   signal load_water_on      : STD_LOGIC;

   signal roura_water_lr     : STD_LOGIC;
   signal roura_water_rl     : STD_LOGIC;
   signal roura_water_bt     : STD_LOGIC;
   signal roura_water_tb     : STD_LOGIC;

   signal roura_water_h        : STD_LOGIC;
   signal roura_water_v        : STD_LOGIC;
   signal roura_water_lenght_1 : unsigned(9 downto 0);
   signal roura_water_lenght_2 : unsigned(9 downto 0);
   signal roura_water_lenght_h : unsigned(9 downto 0);
   signal roura_water_lenght_v : unsigned(9 downto 0);
   signal mini_water_lenght    : unsigned(9 downto 0);
   signal first_water_lenght   : unsigned(9 downto 0);
   signal last_water_lenght    : unsigned(9 downto 0);
   signal roura_water_h_offset : unsigned(9 downto 0);
   signal roura_water_v_offset : unsigned(9 downto 0);

   type rom_type is array (0 to 511) of STD_LOGIC_VECTOR(0 to 31);
   constant ROM : rom_type :=
   (
      "11111111111111111111111111111111",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "10000000000000000000000000000001",
      "11111111111111111111111111111111",

      -- Dalsi obrazek (rovna 1=modra) -- 0001

      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "11100000000000000000000000000111",
      "11100000000000000000000000000111",
      "11100000000000000000000000000111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11100000000000000000000000000111",
      "11100000000000000000000000000111",
      "11100000000000000000000000000111",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",

      -- Dalsi obrazek (zahnuta 1=modra) 0010

      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "11100000000000000000000000000000",
      "11100000000000000000000000000000",
      "11100000000000000000000000000000",
      "11111111111111111111111110000000",
      "11111111111111111111111110000000",
      "11111111111111111111111110000000",
      "11111111111111111111111110000000",
      "11111111111111111111111110000000",
      "11111111111111111111111110000000",
      "11111111111111111111111110000000",
      "00000000000000001111111110000000",
      "00000000000000001111111110000000",
      "00000000000000000011111110000000",
      "00000000000000000011111110000000",
      "11111111111111000011111110000000",
      "11111111111111000011111110000000",
      "11111111111111000011111110000000",
      "11111111111111000011111110000000",
      "11111111111111000011111110000000",
      "11111111111111000011111110000000",
      "11111111111111000011111110000000",
      "11100001111111000011111110000000",
      "11100001111111000011111110000000",
      "11100001111111000011111110000000",
      "00000001111111000011111110000000",
      "00001111111111000011111111110000",
      "00001111111111000011111111110000",
      "00001111111111000011111111110000",

      -- Dalsi obrazek (T 1=modra) - 0011

      "00001111111111000011111111110000",
      "00001111111111000011111111110000",
      "00001111111111000011111111110000",
      "00000001111111000011111110000000",
      "11100001111111000011111110000111",
      "11100001111111000011111110000111",
      "11100001111111000011111110000111",
      "11111111111111000011111111111111",
      "11111111111111000011111111111111",
      "11111111111111000011111111111111",
      "11111111111111000011111111111111",
      "11111111111111000011111111111111",
      "11111111111111000011111111111111",
      "11111111111111000011111111111111",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "11111111111111000011111111111111",
      "11111111111111000011111111111111",
      "11111111111111000011111111111111",
      "11111111111111000011111111111111",
      "11111111111111000011111111111111",
      "11111111111111000011111111111111",
      "11111111111111000011111111111111",
      "11100001111111000011111110000111",
      "11100001111111000011111110000111",
      "11100001111111000011111110000111",
      "00000001111111000011111110000000",
      "00001111111111000011111111110000",
      "00001111111111000011111111110000",
      "00001111111111000011111111110000",

      -- Dalsi obrazek (spodni cast bocni trubky 1=modra) - 0100

      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111001110011100111001110011111",
      "11111001110011100111001110011111",
      "01111111111111111111111111111110",
      "01111111111111111111111111111110",
      "01111111111111111111111111111110",
      "00111111111111111111111111111100",
      "00111111111111111111111111111100",
      "00011111111111111111111111111000",
      "00001111111111111111111111110000",
      "00000111111111111111111111100000",
      "00000011111111111111111111000000",
      "00000001111111111111111110000000",
      "00000000011111111111111000000000",
      "00000000000011111111000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",

      -- Dalsi obrazek (telo trubky 1=bila 8x) - 0101

      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",
      "00100000000000000000000000000100",


      -- Dalsi obrazek (vrchni cast bocni trubky 1=modra) - 0110

      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",

      -- Dalsi obrazek (propojka bocni trubky s hernim polem 1=modra) - 0111

      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "11100000000000000000000000000111",
      "11100000000000000000000000000111",
      "11100000000000000000000000000111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11100000000000000000000000000111",
      "11100000000000000000000000000111",
      "11100000000000000000000000000111",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",

      -- Dalsi obrazek (koncova trubka 1=modra) - 1000

      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "11100000000000000000000000000111",
      "11100000000000000000000000000111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111000011111111111111",
      "11111111111100111100111111111111",
      "11111111111001111110011111111111",
      "11111111111010111101011111111111",
      "11111111110111011011101111111111",
      "11111111110111100111101111111111",
      "11111111110111100111101111111111",
      "11111111110111011011101111111111",
      "11111111111010111101011111111111",
      "11111111111001111110011111111111",
      "11111111111100111100111111111111",
      "11111111111111000011111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11100000000000000000000000000111",
      "11100000000000000000000000000111",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",

      -- text1 (bila) - 1001

      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00011110000111100001111110000111",
      "00011110000111100001111110000111",
      "00011001100110011001100000011000",
      "00011001100110011001100000011000",
      "00011110000111100001111000000110",
      "00011110000111100001111000000110",
      "00011000000110011001100000000001",
      "00011000000110011001100000000001",
      "00011000000110011001111110011110",
      "00011000000110011001111110011110",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000001100001",
      "00000000000000000000000001100001",
      "00000000000000000000000110011001",
      "00000000000000000000000110011001",
      "00000000000000000000000110011001",
      "00000000000000000000000110011001",
      "00000000000000000000000110011001",
      "00000000000000000000000110011001",
      "00000000000000000000000001100001",
      "00000000000000000000000001100001",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",

      -- Dalsi obrazek (tenka trubka ke startovni ohnuta 1=modra) - 1010

      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000000111100000000000000",
      "00000000000001111100000000000000",
      "00000000000011111100000000000000",
      "11111111111111111000000000000000",
      "11111111111111111000000000000000",
      "11111111111111110000000000000000",
      "11111111111111000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",

      -- Dalsi obrazek (tenka trubka ke startovni rovna 1=modra) - 1011

      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "11111111111111111111111111111111",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",

      -- Dalsi obrazek (cihla 1=cervena) - 1100

      "01111111011111110111111101111111",
      "01111111011111110111111101111111",
      "01111111011111110111111101111111",
      "00000000000000000000000000000000",
      "11110111111101111111011111110111",
      "11110111111101111111011111110111",
      "11110111111101111111011111110111",
      "00000000000000000000000000000000",
      "01111111011111110111111101111111",
      "01111111011111110111111101111111",
      "01111111011111110111111101111111",
      "00000000000000000000000000000000",
      "11110111111101111111011111110111",
      "11110111111101111111011111110111",
      "11110111111101111111011111110111",
      "00000000000000000000000000000000",
      "01111111011111110111111101111111",
      "01111111011111110111111101111111",
      "01111111011111110111111101111111",
      "00000000000000000000000000000000",
      "11110111111101111111011111110111",
      "11110111111101111111011111110111",
      "11110111111101111111011111110111",
      "00000000000000000000000000000000",
      "01111111011111110111111101111111",
      "01111111011111110111111101111111",
      "01111111011111110111111101111111",
      "00000000000000000000000000000000",
      "11110111111101111111011111110111",
      "11110111111101111111011111110111",
      "11110111111101111111011111110111",
      "00000000000000000000000000000000",

      -- text2 (bila) - 1101

      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000011000000000011000",
      "00000000000000011000000000011000",
      "10000111100000011000011110011000",
      "10000111100000011000011110011000",
      "00011000000000000001100000000000",
      "00011000000000000001100000000000",
      "00000110000000000000011000000000",
      "00000110000000000000011000000000",
      "10000001100000000000000110000000",
      "10000001100000000000000110000000",
      "00011110000000000001111000000000",
      "00011110000000000001111000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "11100001100110011000011000011001",
      "11100001100110011000011000011001",
      "10011001100110011001100110011001",
      "10011001100110011001100110011001",
      "11100001100110011001100110011001",
      "11100001100110011001100110011001",
      "10011000011000011001100110011001",
      "10011000011000011001100110011001",
      "11100000011000011000011000000110",
      "11100000011000011000011000000110",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",

      -- text3 (bila) - 1110

      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00011111100001100000000001111001",
      "00011111100001100000000001111001",
      "00000110000110011000000110000000",
      "00000110000110011000000110000000",
      "00000110000110011000000001100000",
      "00000110000110011000000001100000",
      "00000110000110011000000000011000",
      "00000110000110011000000000011000",
      "00000110000001100000000111100000",
      "00000110000001100000000111100000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000111100110000001100110000000",
      "00000111100110000001100110000000",
      "00011000000110000001100110000000",
      "00011000000110000001100110000000",
      "00000110000110000000011000000000",
      "00000110000110000000011000000000",
      "00000001100110000000011000000000",
      "00000001100110000000011000000000",
      "00011110000111111000011000011000",
      "00011110000111111000011000011000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",

      -- text4 (bila) - 1111

      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "11111000011000011110000111111000",
      "11111000011000011110000111111000",
      "01100001100110011001100001100000",
      "01100001100110011001100001100000",
      "01100001100110011110000001100000",
      "01100001100110011110000001100000",
      "01100001111110011001100001100000",
      "01100001111110011001100001100000",
      "01100001100110011001100001100000",
      "01100001100110011001100001100000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00011000000000000000000000000000",
      "00011000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",
      "00000000000000000000000000000000",

      others => (others => '0')
   );
   
begin

   pix_x2 <= unsigned(PIXEL_X2);
   pix_y2 <= unsigned(PIXEL_Y2);  

   process (CLK)
   begin
     if rising_edge(CLK) then
         pix_x <= pix_x2;
         pix_y <= pix_y2;
         sig_kurzor  <= KURZOR;
         sig_typ_roury2 <= sig_typ_roury;
      end if;
   end process; 
         sig_komp_on <= KOMP_ON;
         sig_komp_in <= KOMP_IN;

   -- Nastaveni X souradnic pro okraje
   process (CLK) 
   begin
      if (rising_edge(CLK)) then
         if (RST = '1') then
            cell_x_l <= (others => '0');
            cell_x_r <= (others => '0');
         elsif (PIXEL_SET_X = '1' AND GAME_ON = '1') then
            cell_x_l <= pix_x;
            cell_x_r <= pix_x + 31;
         elsif (KOMP_SET_X = '1' AND KOMP_ON = '1') then
            cell_x_l <= pix_x;
            cell_x_r <= pix_x + 31;
         end if;
      end if;
   end process;

   -- Nastaveni Y souradnic pro okraje
   process (CLK) 
   begin
      if (rising_edge(CLK)) then
         if (RST = '1') then
            cell_y_t <= (others => '0');
            cell_y_b <= (others => '0');
         elsif (PIXEL_SET_Y = '1' AND GAME_ON = '1') then
            cell_y_t <= pix_y;
            cell_y_b <= pix_y + 31;
         elsif (KOMP_SET_Y = '1' AND KOMP_ON = '1') then
            cell_y_t <= pix_y;
            cell_y_b <= pix_y + 31;
         end if;
      end if;
   end process;

   -- volba natoceni roury
   sig_natoceni_roury <= sig_komp_in(5 downto 4) when (KOMP_ON = '1')
                      else NATOCENI_ROURY;

   -- volba typu roury
   sig_typ_roury <= sig_komp_in(3 downto 0) when (KOMP_ON = '1')
                    else TYP_ROURY;

   -- Pripraveni souradnic obrazku, rorace obrazku
   process (sig_natoceni_roury, pix_x, pix_y, cell_y_t, cell_x_l)
   begin
      if (sig_natoceni_roury = "01") then -- zahnuta zleva nahoru 01
         img_col  <= 31 - (pix_y(4 downto 0) - cell_y_t(4 downto 0));
         img_row  <= 31 - (pix_x(4 downto 0) - cell_x_l(4 downto 0));
      elsif (sig_natoceni_roury = "10") then -- zahnuta zprava nahoru 10
         img_row  <= 31 - (pix_y(4 downto 0) - cell_y_t(4 downto 0));
         img_col  <= pix_x(4 downto 0) - cell_x_l(4 downto 0);
      elsif (sig_natoceni_roury = "11") then -- zahnuta zprava dolu 11
         img_row  <= pix_y(4 downto 0) - cell_y_t(4 downto 0);
         img_col  <= pix_x(4 downto 0) - cell_x_l(4 downto 0);
      else -- zahnuta zleva dolu 00
         img_row  <= pix_y(4 downto 0) - cell_y_t(4 downto 0);
         img_col  <= 31 - (pix_x(4 downto 0) - cell_x_l(4 downto 0));
      end if;
   end process;

   -- Nastaveni cteci pameti
   rom_addr <= unsigned(sig_typ_roury) & img_row;

   -- Vycteni dat z pameti ROM
   process (CLK)
   begin
      if rising_edge(CLK) then
         rom_data <= ROM(to_integer(rom_addr));  
      end if;
   end process;

   -- Vyber konkretniho bitu ve vyctenem radku obrazku
   rom_bit <= rom_data(to_integer(img_col));

   -- Rika nam ze vykreslujeme pixeli, ktere se nachazi v policku
   sq_cell_on <= '1' when (cell_x_l<=pix_x) and (pix_x<=cell_x_r) and (cell_y_t<=pix_y) and (pix_y<=cell_y_b)
                     else '0';

   --------------------------------------------------------------------
   -- ZOBRAZOVANI VODY V BOCNI ODPOCITAVACI TRUBCE
   --------------------------------------------------------------------

   load_water_lenght <= "00" & (unsigned(LOAD_WATER));

   -- vykresleni vody ktera odpocitava kontrolu trubek
   load_water_on <= '1' when (35 <= pix_x) and (pix_x <= 60) and ((319 - load_water_lenght) <= pix_y) and (pix_y <= 319)
                     else '0';

   --------------------------------------------------------------------
   -- ZOBRAZOVANI VODY V TRUBKACH
   --------------------------------------------------------------------

   process (ZDROJ_VODY1, sig_typ_roury2, ROURA_VODA1, roura_water_lr, roura_water_rl, roura_water_lenght_1, first_water_lenght, last_water_lenght)
   begin
      if ((sig_typ_roury2 = "0001" OR sig_typ_roury2 = "0011") AND ROURA_VODA1(0) = '1' AND ZDROJ_VODY1 = "0001") then
         roura_water_h <= roura_water_lr;
         roura_water_lenght_h <= roura_water_lenght_1;
         roura_water_h_offset <= to_unsigned(0, 10);
      elsif ((sig_typ_roury2 = "0001" OR sig_typ_roury2 = "0011") AND ROURA_VODA1(0) = '1' AND ZDROJ_VODY1 = "0010") then
         roura_water_h <= roura_water_rl;
         roura_water_lenght_h <= roura_water_lenght_1;
         roura_water_h_offset <= to_unsigned(0, 10);
      elsif (sig_typ_roury2 = "0010" AND ROURA_VODA1(0) = '1' AND (ZDROJ_VODY1 = "0101" OR ZDROJ_VODY1 = "0110")) then
         roura_water_h <= roura_water_lr;
         roura_water_lenght_h <= first_water_lenght;
         roura_water_h_offset <= to_unsigned(0, 10);
      elsif (sig_typ_roury2 = "0010" AND ROURA_VODA1(0) = '1' AND (ZDROJ_VODY1 = "0111" OR ZDROJ_VODY1 = "1000")) then
         roura_water_h <= roura_water_rl;
         roura_water_lenght_h <= first_water_lenght;
         roura_water_h_offset <= to_unsigned(0, 10);
      elsif (sig_typ_roury2 = "0010" AND ROURA_VODA1(0) = '1' AND ROURA_VODA1(5) = '1' AND (ZDROJ_VODY1 = "1001" OR ZDROJ_VODY1 = "1011")) then
         roura_water_h <= roura_water_lr;
         roura_water_lenght_h <= last_water_lenght;
         roura_water_h_offset <= to_unsigned(16, 10);
      elsif (sig_typ_roury2 = "0010" AND ROURA_VODA1(0) = '1' AND ROURA_VODA1(5) = '1' AND (ZDROJ_VODY1 = "1010" OR ZDROJ_VODY1 = "1100")) then
         roura_water_h <= roura_water_rl;
         roura_water_lenght_h <= last_water_lenght;
         roura_water_h_offset <= to_unsigned(16, 10);
      else
         roura_water_h <= '0';
         roura_water_lenght_h <= roura_water_lenght_1;
         roura_water_h_offset <= to_unsigned(0, 10);
      end if;
   end process;

   process (ZDROJ_VODY1, ZDROJ_VODY2, sig_typ_roury2, ROURA_VODA1, ROURA_VODA2, roura_water_tb, roura_water_bt,
            roura_water_lenght_2, first_water_lenght, last_water_lenght)
   begin
      if ((sig_typ_roury2 = "0001" OR sig_typ_roury2 = "0011") AND ROURA_VODA2(0) = '1' AND ZDROJ_VODY2 = "0011") then
         roura_water_v <= roura_water_bt;
         roura_water_lenght_v <= roura_water_lenght_2;
         roura_water_v_offset <= to_unsigned(0, 10);
      elsif ((sig_typ_roury2 = "0001" OR sig_typ_roury2 = "0011") AND ROURA_VODA2(0) = '1' AND ZDROJ_VODY2 = "0100") then
         roura_water_v <= roura_water_tb;
         roura_water_lenght_v <= roura_water_lenght_2;
         roura_water_v_offset <= to_unsigned(0, 10);
      elsif (sig_typ_roury2 = "0010" AND ROURA_VODA1(0) = '1' AND ROURA_VODA1(5) = '1' AND (ZDROJ_VODY1 = "0101" OR ZDROJ_VODY1 = "0111")) then
         roura_water_v <= roura_water_bt;
         roura_water_lenght_v <= last_water_lenght;
         roura_water_v_offset <= to_unsigned(16, 10);
      elsif (sig_typ_roury2 = "0010" AND ROURA_VODA1(0) = '1' AND ROURA_VODA1(5) = '1' AND (ZDROJ_VODY1 = "0110" OR ZDROJ_VODY1 = "1000")) then
         roura_water_v <= roura_water_tb;
         roura_water_lenght_v <= last_water_lenght;
         roura_water_v_offset <= to_unsigned(16, 10);
      elsif (sig_typ_roury2 = "0010" AND ROURA_VODA1(0) = '1' AND (ZDROJ_VODY1 = "1010" OR ZDROJ_VODY1 = "1001")) then
         roura_water_v <= roura_water_bt;
         roura_water_lenght_v <= first_water_lenght;
         roura_water_v_offset <= to_unsigned(0, 10);
      elsif (sig_typ_roury2 = "0010" AND ROURA_VODA1(0) = '1' AND (ZDROJ_VODY1 = "1011" OR ZDROJ_VODY1 = "1100")) then
         roura_water_v <= roura_water_tb;
         roura_water_lenght_v <= first_water_lenght;
         roura_water_v_offset <= to_unsigned(0, 10);
      else
         roura_water_v <= '0';
         roura_water_lenght_v <= roura_water_lenght_2;
         roura_water_v_offset <= to_unsigned(0, 10);
      end if;
   end process;

   process (ROURA_VODA1, mini_water_lenght)
   begin
      if (ROURA_VODA1(5) = '1') then
         first_water_lenght <= "0000001111";
         last_water_lenght  <= mini_water_lenght;
      else
         first_water_lenght <= mini_water_lenght;
         last_water_lenght  <= "0000000000";
      end if;
   end process;

   roura_water_lenght_1 <= "00000" & (unsigned(ROURA_VODA1(5 downto 1)));
   roura_water_lenght_2 <= "00000" & (unsigned(ROURA_VODA2(5 downto 1)));
   mini_water_lenght    <= "000000" & (unsigned(ROURA_VODA1(4 downto 1)));
   --------------------------------------------------

   -- zleva doprava 
   roura_water_lr <= '1' when ((cell_x_l + roura_water_h_offset) <= pix_x) and (pix_x <= (cell_x_l + roura_water_h_offset + roura_water_lenght_h))
                        and ((cell_y_t + 14) <= pix_y) and (pix_y <= (cell_y_t + 17))
                     else '0';

   -- zprava doleva
   roura_water_rl <= '1' when (((cell_x_r - roura_water_h_offset) - roura_water_lenght_h) <= pix_x) and (pix_x <= (cell_x_r - roura_water_h_offset))
                        and ((cell_y_t + 14) <= pix_y) and (pix_y <= (cell_y_t + 17))
                     else '0';

   -- zdola nahoru
   roura_water_bt <= '1' when ((cell_x_l + 14) <= pix_x) and (pix_x <= (cell_x_l + 17))
                        and (((cell_y_b - roura_water_v_offset) - roura_water_lenght_v) <= pix_y) and (pix_y <= (cell_y_b - roura_water_v_offset))
                     else '0';

   -- zprava doleva
   roura_water_tb <= '1' when ((cell_x_l + 14) <= pix_x) and (pix_x <= (cell_x_l + 17))
                        and ((cell_y_t + roura_water_v_offset) <= pix_y) and (pix_y <= (cell_y_t + roura_water_v_offset + roura_water_lenght_v))
                     else '0';

   --------------------------------------------------------------------
   -- RIZENI SIGNALU RBG
   --------------------------------------------------------------------

   -- Nastaveni zobrazovane barvy
   process (sq_cell_on, rom_bit, sig_kurzor, sig_typ_roury2, sig_komp_on, pix_x, pix_y, load_water_on, GAME_ON, roura_water_h, roura_water_v)
   begin
      if ((pix_x = 0 AND pix_y = 0) OR (pix_x = 0 AND pix_y = 478) OR (pix_x = 638 AND pix_y = 0) OR (pix_x = 639 AND pix_y = 479)) then
         RGB <= "111";
      elsif (load_water_on = '1' AND GAME_ON = '1') then
         RGB <= "011"; -- voda nacitani
      elsif (roura_water_h = '1' AND sq_cell_on = '1' AND GAME_ON = '1' AND sig_komp_on = '0') then
         RGB <= "011"; -- voda roura nevertikalni
      elsif (roura_water_v = '1' AND sq_cell_on = '1' AND GAME_ON = '1' AND sig_komp_on = '0') then
         RGB <= "011"; -- voda roura vertikalni
      elsif (sq_cell_on = '1' AND rom_bit = '1') then
         if (sig_kurzor = '1' AND sig_komp_on = '0') then
            RGB <= "101";
         elsif (sig_typ_roury2 = "0000" OR sig_typ_roury2 = "1001" OR sig_typ_roury2 = "1101" OR sig_typ_roury2 = "1110" OR sig_typ_roury2 = "1111") then
            RGB <= "111";
         elsif (sig_typ_roury2 = "1100") then
            RGB <= "100";
         else
            RGB <= "001";
         end if;
      else
         RGB <= "000"; 
      end if;
   end process;   

end FULL;